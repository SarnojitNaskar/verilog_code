module NOT_dig(
    input a,
    output b
    );
    assign b=~a;
endmodule
