module comparator_4b_tb;

reg A1, A0, B1, B0;
wire F1, F2, F3;

comparator_4b_dig uut (.A1(A1), .A0(A0), .B1(B1), .B0(B0), .F1(F1), .F2(F2), .F3(F3));

initial
begin
    A1=0;A0=0;B1=0;B0=0;#100;
    A1=0;A0=0;B1=0;B0=1;#100;
    A1=0;A0=0;B1=1;B0=0;#100;
    A1=0;A0=0;B1=1;B0=1;#100;
    A1=0;A0=1;B1=0;B0=0;#100;
    A1=0;A0=1;B1=0;B0=1;#100;
    A1=0;A0=1;B1=1;B0=0;#100;
    A1=0;A0=1;B1=1;B0=1;#100;
    A1=1;A0=0;B1=0;B0=0;#100;
    A1=1;A0=0;B1=0;B0=1;#100;
    A1=1;A0=0;B1=1;B0=0;#100;
    A1=1;A0=0;B1=1;B0=1;#100;
    A1=1;A0=1;B1=0;B0=0;#100;
    A1=1;A0=1;B1=0;B0=1;#100;
    A1=1;A0=1;B1=1;B0=0;#100;
    A1=1;A0=1;B1=1;B0=1;#100;
end
endmodule
