module MUX_41_tb;

reg s1, s0, d0, d1, d2, d3;
wire y;

MUX_41_dig uut (.s1(s1), .s0(s0), .d0(d0), .d1(d1), .d2(d2), .d3(d3), .y(y));

initial
begin
    s1=0;s0=0;d0=1;d1=0;d2=0;d3=0;#100;
    s1=0;s0=0;d0=0;d1=1;d2=1;d3=1;#100;
    s1=0;s0=1;d0=0;d1=1;d2=0;d3=0;#100;
    s1=0;s0=1;d0=1;d1=0;d2=1;d3=1;#100;
    s1=1;s0=0;d0=0;d1=0;d2=1;d3=0;#100;
    s1=1;s0=0;d0=1;d1=1;d2=0;d3=1;#100;
    s1=1;s0=1;d0=0;d1=0;d2=0;d3=1;#100;
    s1=1;s0=1;d0=1;d1=1;d2=1;d3=0;#100;
end

endmodule
