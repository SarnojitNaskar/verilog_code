module mux81_tb;

reg s2, s1, s0;
reg d0, d1, d2, d3, d4, d5, d6, d7;
wire y;

mux_dig uut (.s2(s2), .s1(s1), .s0(s0), 
                .d0(d0), .d1(d1), .d2(d2), .d3(d3), .d4(d4), .d5(d5), .d6(d6), .d7(d7),
                .y(y));

initial
begin
    s2=0;s1=0;s0=0;d0=1;d1=0;d2=0;d3=0;d4=0;d5=0;d6=0;d7=0;#100;
    s2=0;s1=0;s0=0;d0=0;d1=1;d2=1;d3=1;d4=1;d5=1;d6=1;d7=1;#100;
    s2=0;s1=0;s0=1;d0=0;d1=1;d2=0;d3=0;d4=0;d5=0;d6=0;d7=0;#100;
    s2=0;s1=0;s0=1;d0=1;d1=0;d2=1;d3=1;d4=1;d5=1;d6=1;d7=1;#100;
    s2=0;s1=1;s0=0;d0=0;d1=0;d2=1;d3=0;d4=0;d5=0;d6=0;d7=0;#100;
    s2=0;s1=1;s0=0;d0=1;d1=1;d2=0;d3=1;d4=1;d5=1;d6=1;d7=1;#100;
    s2=0;s1=1;s0=1;d0=0;d1=0;d2=0;d3=1;d4=0;d5=0;d6=0;d7=0;#100;
    s2=0;s1=1;s0=1;d0=1;d1=1;d2=1;d3=0;d4=1;d5=1;d6=1;d7=1;#100;
    s2=1;s1=0;s0=0;d0=0;d1=0;d2=0;d3=0;d4=1;d5=0;d6=0;d7=0;#100;
    s2=1;s1=0;s0=0;d0=1;d1=1;d2=1;d3=1;d4=0;d5=1;d6=1;d7=1;#100;
    s2=1;s1=0;s0=1;d0=0;d1=0;d2=0;d3=0;d4=0;d5=1;d6=0;d7=0;#100;
    s2=1;s1=0;s0=1;d0=1;d1=1;d2=1;d3=1;d4=1;d5=0;d6=1;d7=1;#100;
    s2=1;s1=1;s0=0;d0=0;d1=0;d2=0;d3=0;d4=0;d5=0;d6=1;d7=0;#100;
    s2=1;s1=1;s0=0;d0=1;d1=1;d2=1;d3=1;d4=1;d5=1;d6=0;d7=1;#100;
    s2=1;s1=1;s0=1;d0=0;d1=0;d2=0;d3=0;d4=0;d5=0;d6=0;d7=1;#100;
    s2=1;s1=1;s0=1;d0=1;d1=1;d2=1;d3=1;d4=1;d5=1;d6=1;d7=0;#100;
end
endmodule
