module OR_dig(
    input a,
    input b,
    output c
    );
    assign c=a|b;
endmodule
