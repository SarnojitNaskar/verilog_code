module mc_tb;

reg a, b, c;
wire y;

mc_dig uut (.a(a), .b(b), .c(c), .y(y));

initial
begin
    a=0;b=0;c=0;#100;
    a=0;b=0;c=1;#100;
    a=0;b=1;c=0;#100;
    a=0;b=1;c=1;#100;
    a=1;b=0;c=0;#100;
    a=1;b=0;c=1;#100;
    a=1;b=1;c=0;#100;
    a=1;b=1;c=1;#100;
end
endmodule
